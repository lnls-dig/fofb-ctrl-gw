`define WB_FOFB_PROCESSING_REGS_SIZE 26624
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_FIXED_POINT_POS 'h0
`define WB_FOFB_PROCESSING_REGS_COEFFS_FIXED_POINT_POS_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_COEFFS_FIXED_POINT_POS_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_0 'h800
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_0_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_0_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_1 'h1000
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_1_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_1_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_2 'h1800
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_2_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_2_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_3 'h2000
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_3_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_3_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_4 'h2800
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_4_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_4_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_5 'h3000
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_5_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_5_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_6 'h3800
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_6_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_6_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_7 'h4000
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_7_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_7_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_8 'h4800
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_8_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_8_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_9 'h5000
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_9_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_9_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_10 'h5800
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_10_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_10_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_11 'h6000
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_11_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_11_DATA 'h0
