`define WB_FOFB_PROCESSING_REGS_SIZE 12
`define ADDR_WB_FOFB_PROCESSING_REGS_RAM_COEFF_DAT 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_RAM_COEFF_ADDR 'h4
`define ADDR_WB_FOFB_PROCESSING_REGS_RAM_WRITE 'h8
`define WB_FOFB_PROCESSING_REGS_RAM_WRITE_ENABLE_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_RAM_WRITE_ENABLE 'h1
