`define WB_FOFB_PROCESSING_REGS_SIZE 16
`define ADDR_WB_FOFB_PROCESSING_REGS_RAM_WRITE 'h0
`define WB_FOFB_PROCESSING_REGS_RAM_WRITE_ENABLE_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_RAM_WRITE_ENABLE 'h1
`define ADDR_WB_FOFB_PROCESSING_REGS_RAM_DATA_IN 'h4
`define WB_FOFB_PROCESSING_REGS_RAM_DATA_IN_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_RAM_DATA_IN_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_RAM_DATA_OUT 'h8
`define WB_FOFB_PROCESSING_REGS_RAM_DATA_OUT_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_RAM_DATA_OUT_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_RAM_ADDR 'hc
`define WB_FOFB_PROCESSING_REGS_RAM_ADDR_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_RAM_ADDR_VAL 'hfff
