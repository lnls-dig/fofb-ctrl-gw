package wb_fofb_processing_regs_consts_pkg is
  constant c_WB_FOFB_PROCESSING_REGS_SIZE : Natural := 28672;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_FIXED_POINT_POS_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_FIXED_POINT_POS_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACCS_GAINS_FIXED_POINT_POS_ADDR : Natural := 16#4#;
  constant c_WB_FOFB_PROCESSING_REGS_ACCS_GAINS_FIXED_POINT_POS_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_0_ADDR : Natural := 16#8#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_0_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_0_ADDR : Natural := 16#c#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_0_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_0_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_1_ADDR : Natural := 16#10#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_1_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_1_ADDR : Natural := 16#14#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_1_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_1_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_2_ADDR : Natural := 16#18#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_2_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_2_ADDR : Natural := 16#1c#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_2_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_2_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_3_ADDR : Natural := 16#20#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_3_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_3_ADDR : Natural := 16#24#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_3_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_3_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_4_ADDR : Natural := 16#28#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_4_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_4_ADDR : Natural := 16#2c#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_4_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_4_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_5_ADDR : Natural := 16#30#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_5_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_5_ADDR : Natural := 16#34#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_5_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_5_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_6_ADDR : Natural := 16#38#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_6_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_6_ADDR : Natural := 16#3c#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_6_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_6_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_7_ADDR : Natural := 16#40#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_7_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_7_ADDR : Natural := 16#44#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_7_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_7_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_8_ADDR : Natural := 16#48#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_8_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_8_ADDR : Natural := 16#4c#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_8_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_8_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_9_ADDR : Natural := 16#50#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_9_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_9_ADDR : Natural := 16#54#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_9_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_9_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_10_ADDR : Natural := 16#58#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_10_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_10_ADDR : Natural := 16#5c#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_10_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_10_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_11_ADDR : Natural := 16#60#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_GAIN_11_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_11_ADDR : Natural := 16#64#;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_11_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_ACC_CTL_11_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_0_ADDR : Natural := 16#68#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_0_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_0_ADDR : Natural := 16#6c#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_0_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_1_ADDR : Natural := 16#70#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_1_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_1_ADDR : Natural := 16#74#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_1_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_2_ADDR : Natural := 16#78#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_2_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_2_ADDR : Natural := 16#7c#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_2_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_3_ADDR : Natural := 16#80#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_3_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_3_ADDR : Natural := 16#84#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_3_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_4_ADDR : Natural := 16#88#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_4_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_4_ADDR : Natural := 16#8c#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_4_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_5_ADDR : Natural := 16#90#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_5_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_5_ADDR : Natural := 16#94#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_5_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_6_ADDR : Natural := 16#98#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_6_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_6_ADDR : Natural := 16#9c#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_6_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_7_ADDR : Natural := 16#a0#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_7_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_7_ADDR : Natural := 16#a4#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_7_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_8_ADDR : Natural := 16#a8#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_8_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_8_ADDR : Natural := 16#ac#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_8_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_9_ADDR : Natural := 16#b0#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_9_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_9_ADDR : Natural := 16#b4#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_9_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_10_ADDR : Natural := 16#b8#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_10_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_10_ADDR : Natural := 16#bc#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_10_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_11_ADDR : Natural := 16#c0#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MAX_11_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_11_ADDR : Natural := 16#c4#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_MIN_11_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_0_ADDR : Natural := 16#800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_0_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_0_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_1_ADDR : Natural := 16#1000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_1_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_1_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_2_ADDR : Natural := 16#1800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_2_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_2_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_3_ADDR : Natural := 16#2000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_3_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_3_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_4_ADDR : Natural := 16#2800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_4_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_4_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_5_ADDR : Natural := 16#3000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_5_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_5_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_6_ADDR : Natural := 16#3800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_6_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_6_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_7_ADDR : Natural := 16#4000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_7_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_7_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_8_ADDR : Natural := 16#4800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_8_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_8_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_9_ADDR : Natural := 16#5000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_9_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_9_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_10_ADDR : Natural := 16#5800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_10_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_10_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_11_ADDR : Natural := 16#6000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_11_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_11_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_SETPOINTS_RAM_BANK_ADDR : Natural := 16#6800#;
  constant c_WB_FOFB_PROCESSING_REGS_SETPOINTS_RAM_BANK_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_SETPOINTS_RAM_BANK_DATA_ADDR : Natural := 16#0#;
end package wb_fofb_processing_regs_consts_pkg;
