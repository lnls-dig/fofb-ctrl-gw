`define FOFB_CC_CSR_SIZE 8196
`define ADDR_FOFB_CC_CSR_RAM_REG 'h0
`define FOFB_CC_CSR_RAM_REG_SIZE 4
`define ADDR_FOFB_CC_CSR_RAM_REG_DATA 'h0
`define ADDR_FOFB_CC_CSR_CFG_VAL 'h2000
