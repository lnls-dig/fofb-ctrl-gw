`define FOFB_CC_CSR_SIZE 16384
`define ADDR_FOFB_CC_CSR_CFG_VAL 'h0
`define ADDR_FOFB_CC_CSR_CFG_CTL 'h4
`define FOFB_CC_CSR_CFG_CTL_READ_RAM_OFFSET 0
`define FOFB_CC_CSR_CFG_CTL_READ_RAM 'h1
`define ADDR_FOFB_CC_CSR_RAM_REG 'h2000
`define FOFB_CC_CSR_RAM_REG_SIZE 4
`define ADDR_FOFB_CC_CSR_RAM_REG_DATA 'h0
