package wb_fofb_sys_id_regs_consts_pkg is
  constant c_WB_FOFB_SYS_ID_REGS_SIZE : Natural := 8;
  constant c_WB_FOFB_SYS_ID_REGS_BPM_POS_FLATENIZER_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_SYS_ID_REGS_BPM_POS_FLATENIZER_SIZE : Natural := 8;
  constant c_WB_FOFB_SYS_ID_REGS_BPM_POS_FLATENIZER_MAX_NUM_CTE_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_SYS_ID_REGS_BPM_POS_FLATENIZER_BASE_BPM_ID_ADDR : Natural := 16#4#;
end package wb_fofb_sys_id_regs_consts_pkg;
