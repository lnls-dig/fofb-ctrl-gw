`define WB_FOFB_PROCESSING_REGS_SIZE 28672
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_FIXED_POINT_POS 'h0
`define WB_FOFB_PROCESSING_REGS_COEFFS_FIXED_POINT_POS_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_COEFFS_FIXED_POINT_POS_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_ACCS_GAINS_FIXED_POINT_POS 'h4
`define WB_FOFB_PROCESSING_REGS_ACCS_GAINS_FIXED_POINT_POS_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACCS_GAINS_FIXED_POINT_POS_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_GAIN_0 'h8
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_0_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_0_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_CTL_0 'hc
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_0_CLEAR_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_0_CLEAR 'h1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_0_FREEZE_OFFSET 1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_0_FREEZE 'h2
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_GAIN_1 'h10
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_1_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_1_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_CTL_1 'h14
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_1_CLEAR_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_1_CLEAR 'h1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_1_FREEZE_OFFSET 1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_1_FREEZE 'h2
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_GAIN_2 'h18
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_2_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_2_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_CTL_2 'h1c
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_2_CLEAR_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_2_CLEAR 'h1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_2_FREEZE_OFFSET 1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_2_FREEZE 'h2
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_GAIN_3 'h20
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_3_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_3_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_CTL_3 'h24
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_3_CLEAR_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_3_CLEAR 'h1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_3_FREEZE_OFFSET 1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_3_FREEZE 'h2
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_GAIN_4 'h28
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_4_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_4_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_CTL_4 'h2c
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_4_CLEAR_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_4_CLEAR 'h1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_4_FREEZE_OFFSET 1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_4_FREEZE 'h2
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_GAIN_5 'h30
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_5_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_5_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_CTL_5 'h34
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_5_CLEAR_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_5_CLEAR 'h1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_5_FREEZE_OFFSET 1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_5_FREEZE 'h2
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_GAIN_6 'h38
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_6_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_6_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_CTL_6 'h3c
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_6_CLEAR_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_6_CLEAR 'h1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_6_FREEZE_OFFSET 1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_6_FREEZE 'h2
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_GAIN_7 'h40
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_7_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_7_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_CTL_7 'h44
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_7_CLEAR_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_7_CLEAR 'h1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_7_FREEZE_OFFSET 1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_7_FREEZE 'h2
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_GAIN_8 'h48
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_8_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_8_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_CTL_8 'h4c
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_8_CLEAR_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_8_CLEAR 'h1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_8_FREEZE_OFFSET 1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_8_FREEZE 'h2
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_GAIN_9 'h50
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_9_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_9_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_CTL_9 'h54
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_9_CLEAR_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_9_CLEAR 'h1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_9_FREEZE_OFFSET 1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_9_FREEZE 'h2
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_GAIN_10 'h58
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_10_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_10_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_CTL_10 'h5c
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_10_CLEAR_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_10_CLEAR 'h1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_10_FREEZE_OFFSET 1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_10_FREEZE 'h2
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_GAIN_11 'h60
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_11_VAL_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_GAIN_11_VAL 'hffffffff
`define ADDR_WB_FOFB_PROCESSING_REGS_ACC_CTL_11 'h64
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_11_CLEAR_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_11_CLEAR 'h1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_11_FREEZE_OFFSET 1
`define WB_FOFB_PROCESSING_REGS_ACC_CTL_11_FREEZE 'h2
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_0 'h800
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_0_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_0_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_1 'h1000
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_1_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_1_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_2 'h1800
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_2_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_2_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_3 'h2000
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_3_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_3_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_4 'h2800
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_4_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_4_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_5 'h3000
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_5_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_5_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_6 'h3800
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_6_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_6_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_7 'h4000
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_7_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_7_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_8 'h4800
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_8_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_8_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_9 'h5000
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_9_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_9_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_10 'h5800
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_10_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_10_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_11 'h6000
`define WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_11_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_11_DATA 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_SETPOINTS_RAM_BANK 'h6800
`define WB_FOFB_PROCESSING_REGS_SETPOINTS_RAM_BANK_SIZE 4
`define ADDR_WB_FOFB_PROCESSING_REGS_SETPOINTS_RAM_BANK_DATA 'h0
