`define WB_FOFB_PROCESSING_REGS_SIZE 16
`define ADDR_WB_FOFB_PROCESSING_REGS_RAM_DATA_IN 'h0
`define ADDR_WB_FOFB_PROCESSING_REGS_RAM_DATA_OUT 'h4
`define ADDR_WB_FOFB_PROCESSING_REGS_RAM_ADDR 'h8
`define ADDR_WB_FOFB_PROCESSING_REGS_RAM_WRITE 'hc
`define WB_FOFB_PROCESSING_REGS_RAM_WRITE_ENABLE_OFFSET 0
`define WB_FOFB_PROCESSING_REGS_RAM_WRITE_ENABLE 'h1
