package wb_fofb_processing_regs_consts_pkg is
  constant c_WB_FOFB_PROCESSING_REGS_SIZE : Natural := 28672;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_FIXED_POINT_POS_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_FIXED_POINT_POS_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_0_ADDR : Natural := 16#800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_0_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_0_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_1_ADDR : Natural := 16#1000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_1_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_1_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_2_ADDR : Natural := 16#1800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_2_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_2_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_3_ADDR : Natural := 16#2000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_3_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_3_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_4_ADDR : Natural := 16#2800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_4_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_4_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_5_ADDR : Natural := 16#3000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_5_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_5_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_6_ADDR : Natural := 16#3800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_6_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_6_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_7_ADDR : Natural := 16#4000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_7_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_7_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_8_ADDR : Natural := 16#4800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_8_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_8_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_9_ADDR : Natural := 16#5000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_9_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_9_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_10_ADDR : Natural := 16#5800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_10_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_10_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_11_ADDR : Natural := 16#6000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_11_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_11_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_SETPOINTS_RAM_BANK_ADDR : Natural := 16#6800#;
  constant c_WB_FOFB_PROCESSING_REGS_SETPOINTS_RAM_BANK_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_SETPOINTS_RAM_BANK_DATA_ADDR : Natural := 16#0#;
end package wb_fofb_processing_regs_consts_pkg;
