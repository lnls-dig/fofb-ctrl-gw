package wb_fofb_processing_regs_consts_pkg is
  constant c_WB_FOFB_PROCESSING_REGS_SIZE : natural := 26624;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_FIXED_POINT_POS : natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_FIXED_POINT_POS_VAL_OFFSET : natural := 0;
--  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_FIXED_POINT_POS_VAL : natural := 16#ffffffff#; NOTE: violates bounds
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_0 : natural := 16#800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_0_SIZE : natural := 4;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_0_DATA : natural := 16#0#;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_1 : natural := 16#1000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_1_SIZE : natural := 4;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_1_DATA : natural := 16#0#;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_2 : natural := 16#1800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_2_SIZE : natural := 4;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_2_DATA : natural := 16#0#;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_3 : natural := 16#2000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_3_SIZE : natural := 4;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_3_DATA : natural := 16#0#;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_4 : natural := 16#2800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_4_SIZE : natural := 4;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_4_DATA : natural := 16#0#;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_5 : natural := 16#3000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_5_SIZE : natural := 4;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_5_DATA : natural := 16#0#;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_6 : natural := 16#3800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_6_SIZE : natural := 4;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_6_DATA : natural := 16#0#;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_7 : natural := 16#4000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_7_SIZE : natural := 4;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_7_DATA : natural := 16#0#;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_8 : natural := 16#4800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_8_SIZE : natural := 4;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_8_DATA : natural := 16#0#;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_9 : natural := 16#5000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_9_SIZE : natural := 4;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_9_DATA : natural := 16#0#;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_10 : natural := 16#5800#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_10_SIZE : natural := 4;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_10_DATA : natural := 16#0#;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_11 : natural := 16#6000#;
  constant c_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_11_SIZE : natural := 4;
  constant c_ADDR_WB_FOFB_PROCESSING_REGS_COEFFS_RAM_BANK_11_DATA : natural := 16#0#;
end package wb_fofb_processing_regs_consts_pkg;
