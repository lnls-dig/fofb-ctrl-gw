`define MATMUL_WB_SIZE 12
`define ADDR_MATMUL_WB_RAM_COEFF_DAT 'h0
`define ADDR_MATMUL_WB_RAM_COEFF_ADDR 'h4
`define ADDR_MATMUL_WB_RAM_WRITE 'h8
`define MATMUL_WB_RAM_WRITE_ENABLE_OFFSET 0
`define MATMUL_WB_RAM_WRITE_ENABLE 'h1
