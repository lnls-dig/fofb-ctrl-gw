`define FOFB_CC_REGS_SIZE 16384
`define ADDR_FOFB_CC_REGS_CFG_VAL 'h0
`define FOFB_CC_REGS_CFG_VAL_ACT_PART_OFFSET 0
`define FOFB_CC_REGS_CFG_VAL_ACT_PART 'h1
`define FOFB_CC_REGS_CFG_VAL_UNUSED_OFFSET 1
`define FOFB_CC_REGS_CFG_VAL_UNUSED 'h2
`define FOFB_CC_REGS_CFG_VAL_ERR_CLR_OFFSET 2
`define FOFB_CC_REGS_CFG_VAL_ERR_CLR 'h4
`define FOFB_CC_REGS_CFG_VAL_CC_ENABLE_OFFSET 3
`define FOFB_CC_REGS_CFG_VAL_CC_ENABLE 'h8
`define FOFB_CC_REGS_CFG_VAL_TFS_OVERRIDE_OFFSET 4
`define FOFB_CC_REGS_CFG_VAL_TFS_OVERRIDE 'h10
`define ADDR_FOFB_CC_REGS_TOA_CTL 'h4
`define FOFB_CC_REGS_TOA_CTL_RD_EN_OFFSET 0
`define FOFB_CC_REGS_TOA_CTL_RD_EN 'h1
`define FOFB_CC_REGS_TOA_CTL_RD_STR_OFFSET 1
`define FOFB_CC_REGS_TOA_CTL_RD_STR 'h2
`define ADDR_FOFB_CC_REGS_TOA_DATA 'h8
`define FOFB_CC_REGS_TOA_DATA_VAL_OFFSET 0
`define FOFB_CC_REGS_TOA_DATA_VAL 'hffffffff
`define ADDR_FOFB_CC_REGS_RCB_CTL 'hc
`define FOFB_CC_REGS_RCB_CTL_RD_EN_OFFSET 0
`define FOFB_CC_REGS_RCB_CTL_RD_EN 'h1
`define FOFB_CC_REGS_RCB_CTL_RD_STR_OFFSET 1
`define FOFB_CC_REGS_RCB_CTL_RD_STR 'h2
`define ADDR_FOFB_CC_REGS_RCB_DATA 'h10
`define FOFB_CC_REGS_RCB_DATA_VAL_OFFSET 0
`define FOFB_CC_REGS_RCB_DATA_VAL 'hffffffff
`define ADDR_FOFB_CC_REGS_RAM_REG 'h2000
`define FOFB_CC_REGS_RAM_REG_SIZE 4
`define ADDR_FOFB_CC_REGS_RAM_REG_DATA 'h0
