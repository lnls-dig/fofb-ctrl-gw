-------------------------------------------------------------------------------
-- Title      :  Dot product package
-------------------------------------------------------------------------------
-- Author     :  Melissa Aguiar
-- Company    :  CNPEM LNLS-DIG
-- Platform   :  FPGA-generic
-------------------------------------------------------------------------------
-- Description:  Package for the dot product core
-------------------------------------------------------------------------------
-- Copyright (c) 2020 CNPEM
-- Licensed under GNU Lesser General Public License (LGPL) v3.0
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author                Description
-- 2021-07-30  1.0      melissa.aguiar        Created
-- 2022-07-27  1.1      guilherme.ricioli     Changed coeffs RAMs' wb interface
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package dot_prod_pkg is

  -- fofb_processing output array
  -- NOTE:  c_Q_WIDTH must match with g_Q_WIDTH defined on
  --        hdl/top/afc_ref_design_gen/afc_ref_fofb_ctrl_gen.vhd
  constant c_Q_WIDTH               : natural := 16;
  type t_fofb_processing_setpoints is array (natural range <>) of signed(c_Q_WIDTH-1 downto 0);

  -- Input record
  type t_dot_prod_record_fod is record
    valid                        : std_logic;
    data                         : std_logic_vector(32-1 downto 0);
    addr                         : std_logic_vector(9-1 downto 0);
  end record t_dot_prod_record_fod;

  -- Input array of record
  type t_dot_prod_array_record_fod is array (natural range <>) of t_dot_prod_record_fod;

  -- RAM interface arrays
  -- NOTE:  These values must agree with c_ADDR_WIDTH and c_DATA_WIDTH defined on
  --        hdl/top/afc_ref_design_gen/afc_ref_fofb_ctrl_gen.vhd
  constant c_ADDR_WIDTH_cp         : natural := 9;
  constant c_DATA_WIDTH_cp         : natural := 32;
  type t_arr_coeff_ram_addr is array (natural range <>) of std_logic_vector(c_ADDR_WIDTH_cp-1 downto 0);
  type t_arr_coeff_ram_data is array (natural range <>) of std_logic_vector(c_DATA_WIDTH_cp-1 downto 0);

  component dot_prod is
    generic(
      -- Width for input a[k]
      g_A_WIDTH                    : natural := 32;

      -- Width for input b[k]
      g_B_WIDTH                    : natural := 32;

      -- Width for output
      g_C_WIDTH                    : natural := 16;

      -- Fixed point representation for output
      g_OUT_FIXED                  : natural := 26;

      -- Extra bits for accumulator
      g_EXTRA_WIDTH                : natural := 4
    );
    port(
      -- Core clock
      clk_i                        : in std_logic;

      -- Reset
      rst_n_i                      : in std_logic;

      -- Clear
      clear_acc_i                  : in std_logic;

      -- Data valid input
      valid_i                      : in std_logic;

      -- Time frame end
      time_frame_end_i             : in std_logic;

      -- Input a[k]
      a_i                          : in signed(g_A_WIDTH-1 downto 0);

      -- Input b[k]
      b_i                          : in signed(g_B_WIDTH-1 downto 0);

      -- Result output
      result_o                     : out signed(g_C_WIDTH-1 downto 0);
      result_debug_o               : out signed(g_C_WIDTH-1 downto 0);

      -- Data valid output
      result_valid_end_o           : out std_logic;
      result_valid_debug_o         : out std_logic
    );
  end component dot_prod;

  component dot_prod_coeff_vec is
    generic(
      -- Width for DCC input
      g_A_WIDTH                    : natural := 32;

      -- Width for DCC addr
      g_ID_WIDTH                   : natural := 9;

      -- Width for RAM coeff
      g_B_WIDTH                    : natural;

      -- Width for RAM addr
      g_K_WIDTH                    : natural;

      -- Width for output
      g_C_WIDTH                    : natural := 16;

      -- Fixed point representation for output
      g_OUT_FIXED                  : natural := 26;

      -- Extra bits for accumulator
      g_EXTRA_WIDTH                : natural := 4
    );
    port(
      -- Core clock
      clk_i                        : in std_logic;

      -- Reset
      rst_n_i                      : in std_logic;

      -- DCC interface
      dcc_valid_i                  : in std_logic;
      dcc_data_i                   : in signed(g_A_WIDTH-1 downto 0);
      dcc_addr_i                   : in std_logic_vector(g_ID_WIDTH-1 downto 0);
      dcc_time_frame_start_i       : in std_logic;
      dcc_time_frame_end_i         : in std_logic;

      -- RAM interface
      coeff_ram_addr_o             : out std_logic_vector(g_K_WIDTH-1 downto 0);
      coeff_ram_data_i             : in std_logic_vector(g_B_WIDTH-1 downto 0);

      -- Result output array
      sp_o                         : out signed(g_C_WIDTH-1 downto 0);
      sp_debug_o                   : out signed(g_C_WIDTH-1 downto 0);

      -- Valid output
      sp_valid_o                   : out std_logic;
      sp_valid_debug_o             : out std_logic
    );
  end component dot_prod_coeff_vec;

  component fofb_processing_channel is
    generic(
      -- Width for DCC input
      g_A_WIDTH                    : natural := 32;

      -- Width for DCC addr
      g_ID_WIDTH                   : natural := 9;

      -- Width for RAM coeff
      g_B_WIDTH                    : natural;

      -- Width for RAM addr
      g_K_WIDTH                    : natural;

      -- Width for output
      g_C_WIDTH                    : natural := 16;

      -- Fixed point representation for output
      g_OUT_FIXED                  : natural := 26;

      -- Extra bits for accumulator
      g_EXTRA_WIDTH                : natural := 4;

      g_ANTI_WINDUP_UPPER_LIMIT    : integer; -- anti-windup upper limit
      g_ANTI_WINDUP_LOWER_LIMIT    : integer  -- anti-windup lower limit
    );
    port(
      ---------------------------------------------------------------------------
      -- Clock and reset interface
      ---------------------------------------------------------------------------
      clk_i                        : in std_logic;
      rst_n_i                      : in std_logic;

      ---------------------------------------------------------------------------
      -- Dot product Interface Signals
      ---------------------------------------------------------------------------
      -- DCC interface
      dcc_valid_i                  : in std_logic;
      dcc_data_i                   : in signed(g_A_WIDTH-1 downto 0);
      dcc_addr_i                   : in std_logic_vector(g_ID_WIDTH-1 downto 0);
      dcc_time_frame_start_i       : in std_logic;
      dcc_time_frame_end_i         : in std_logic;

      -- RAM interface
      coeff_ram_addr_o             : out std_logic_vector(g_K_WIDTH-1 downto 0);
      coeff_ram_data_i             : in std_logic_vector(g_B_WIDTH-1 downto 0);

      -- Setpoint
      sp_o                         : out signed(g_C_WIDTH-1 downto 0);
      sp_valid_o                   : out std_logic
    );
  end component fofb_processing_channel;

  component fofb_processing is
    generic(
      -- Width for DCC input
      g_A_WIDTH                    : natural := 32;

      -- Width for DCC addr
      g_ID_WIDTH                   : natural := 9;

      -- Width for RAM coeff
      g_B_WIDTH                    : natural;

      -- Width for RAM addr
      g_K_WIDTH                    : natural;

      -- Width for output
      g_C_WIDTH                    : natural := 16;

      -- Fixed point representation for output
      g_OUT_FIXED                  : natural := 26;

      -- Extra bits for accumulator
      g_EXTRA_WIDTH                : natural := 4;

      -- Number of channels
      g_CHANNELS                   : natural;

      g_ANTI_WINDUP_UPPER_LIMIT    : integer; -- anti-windup upper limit
      g_ANTI_WINDUP_LOWER_LIMIT    : integer  -- anti-windup lower limit
    );
    port(
      ---------------------------------------------------------------------------
      -- FOFB processing channel interface
      ---------------------------------------------------------------------------
      -- Clock core
      clk_i                        : in std_logic;

      -- Reset
      rst_n_i                      : in std_logic;

      -- DCC interface
      dcc_fod_i                    : in t_dot_prod_array_record_fod;
      dcc_time_frame_start_i       : in std_logic;
      dcc_time_frame_end_i    	   : in std_logic;

      -- RAM interface
      coeff_ram_addr_arr_o         : out t_arr_coeff_ram_addr;
      coeff_ram_data_arr_i         : in t_arr_coeff_ram_data;

      -- Setpoints
      sp_arr_o                     : out t_fofb_processing_setpoints(g_CHANNELS-1 downto 0);
      sp_valid_arr_o               : out std_logic_vector(g_CHANNELS-1 downto 0)
    );
  end component fofb_processing;

  component wb_fofb_processing_regs is
    port (
      rst_n_i              : in    std_logic;
      clk_sys_i            : in    std_logic;
      wb_adr_i             : in    std_logic_vector(12 downto 0);
      wb_dat_i             : in    std_logic_vector(31 downto 0);
      wb_dat_o             : out   std_logic_vector(31 downto 0);
      wb_cyc_i             : in    std_logic;
      wb_sel_i             : in    std_logic_vector(3 downto 0);
      wb_stb_i             : in    std_logic;
      wb_we_i              : in    std_logic;
      wb_ack_o             : out   std_logic;
      wb_stall_o           : out   std_logic;
      wb_fofb_processing_regs_clk_i : in    std_logic;
      -- Ports for RAM: FOFB PROCESSING RAM bank for register map
      wb_fofb_processing_regs_ram_bank_0_addr_i : in    std_logic_vector(8 downto 0);
      -- Read data output
      wb_fofb_processing_regs_ram_bank_0_data_o : out   std_logic_vector(31 downto 0);
      -- Read strobe input (active high)
      wb_fofb_processing_regs_ram_bank_0_rd_i : in    std_logic;
      -- Write data input
      wb_fofb_processing_regs_ram_bank_0_data_i : in    std_logic_vector(31 downto 0);
      -- Write strobe (active high)
      wb_fofb_processing_regs_ram_bank_0_wr_i : in    std_logic;
      -- Ports for RAM: FOFB PROCESSING RAM bank for register map
      wb_fofb_processing_regs_ram_bank_1_addr_i : in    std_logic_vector(8 downto 0);
      -- Read data output
      wb_fofb_processing_regs_ram_bank_1_data_o : out   std_logic_vector(31 downto 0);
      -- Read strobe input (active high)
      wb_fofb_processing_regs_ram_bank_1_rd_i : in    std_logic;
      -- Write data input
      wb_fofb_processing_regs_ram_bank_1_data_i : in    std_logic_vector(31 downto 0);
      -- Write strobe (active high)
      wb_fofb_processing_regs_ram_bank_1_wr_i : in    std_logic;
      -- Ports for RAM: FOFB PROCESSING RAM bank for register map
      wb_fofb_processing_regs_ram_bank_2_addr_i : in    std_logic_vector(8 downto 0);
      -- Read data output
      wb_fofb_processing_regs_ram_bank_2_data_o : out   std_logic_vector(31 downto 0);
      -- Read strobe input (active high)
      wb_fofb_processing_regs_ram_bank_2_rd_i : in    std_logic;
      -- Write data input
      wb_fofb_processing_regs_ram_bank_2_data_i : in    std_logic_vector(31 downto 0);
      -- Write strobe (active high)
      wb_fofb_processing_regs_ram_bank_2_wr_i : in    std_logic;
      -- Ports for RAM: FOFB PROCESSING RAM bank for register map
      wb_fofb_processing_regs_ram_bank_3_addr_i : in    std_logic_vector(8 downto 0);
      -- Read data output
      wb_fofb_processing_regs_ram_bank_3_data_o : out   std_logic_vector(31 downto 0);
      -- Read strobe input (active high)
      wb_fofb_processing_regs_ram_bank_3_rd_i : in    std_logic;
      -- Write data input
      wb_fofb_processing_regs_ram_bank_3_data_i : in    std_logic_vector(31 downto 0);
      -- Write strobe (active high)
      wb_fofb_processing_regs_ram_bank_3_wr_i : in    std_logic;
      -- Ports for RAM: FOFB PROCESSING RAM bank for register map
      wb_fofb_processing_regs_ram_bank_4_addr_i : in    std_logic_vector(8 downto 0);
      -- Read data output
      wb_fofb_processing_regs_ram_bank_4_data_o : out   std_logic_vector(31 downto 0);
      -- Read strobe input (active high)
      wb_fofb_processing_regs_ram_bank_4_rd_i : in    std_logic;
      -- Write data input
      wb_fofb_processing_regs_ram_bank_4_data_i : in    std_logic_vector(31 downto 0);
      -- Write strobe (active high)
      wb_fofb_processing_regs_ram_bank_4_wr_i : in    std_logic;
      -- Ports for RAM: FOFB PROCESSING RAM bank for register map
      wb_fofb_processing_regs_ram_bank_5_addr_i : in    std_logic_vector(8 downto 0);
      -- Read data output
      wb_fofb_processing_regs_ram_bank_5_data_o : out   std_logic_vector(31 downto 0);
      -- Read strobe input (active high)
      wb_fofb_processing_regs_ram_bank_5_rd_i : in    std_logic;
      -- Write data input
      wb_fofb_processing_regs_ram_bank_5_data_i : in    std_logic_vector(31 downto 0);
      -- Write strobe (active high)
      wb_fofb_processing_regs_ram_bank_5_wr_i : in    std_logic;
      -- Ports for RAM: FOFB PROCESSING RAM bank for register map
      wb_fofb_processing_regs_ram_bank_6_addr_i : in    std_logic_vector(8 downto 0);
      -- Read data output
      wb_fofb_processing_regs_ram_bank_6_data_o : out   std_logic_vector(31 downto 0);
      -- Read strobe input (active high)
      wb_fofb_processing_regs_ram_bank_6_rd_i : in    std_logic;
      -- Write data input
      wb_fofb_processing_regs_ram_bank_6_data_i : in    std_logic_vector(31 downto 0);
      -- Write strobe (active high)
      wb_fofb_processing_regs_ram_bank_6_wr_i : in    std_logic;
      -- Ports for RAM: FOFB PROCESSING RAM bank for register map
      wb_fofb_processing_regs_ram_bank_7_addr_i : in    std_logic_vector(8 downto 0);
      -- Read data output
      wb_fofb_processing_regs_ram_bank_7_data_o : out   std_logic_vector(31 downto 0);
      -- Read strobe input (active high)
      wb_fofb_processing_regs_ram_bank_7_rd_i : in    std_logic;
      -- Write data input
      wb_fofb_processing_regs_ram_bank_7_data_i : in    std_logic_vector(31 downto 0);
      -- Write strobe (active high)
      wb_fofb_processing_regs_ram_bank_7_wr_i : in    std_logic;
      -- Ports for RAM: FOFB PROCESSING RAM bank for register map
      wb_fofb_processing_regs_ram_bank_8_addr_i : in    std_logic_vector(8 downto 0);
      -- Read data output
      wb_fofb_processing_regs_ram_bank_8_data_o : out   std_logic_vector(31 downto 0);
      -- Read strobe input (active high)
      wb_fofb_processing_regs_ram_bank_8_rd_i : in    std_logic;
      -- Write data input
      wb_fofb_processing_regs_ram_bank_8_data_i : in    std_logic_vector(31 downto 0);
      -- Write strobe (active high)
      wb_fofb_processing_regs_ram_bank_8_wr_i : in    std_logic;
      -- Ports for RAM: FOFB PROCESSING RAM bank for register map
      wb_fofb_processing_regs_ram_bank_9_addr_i : in    std_logic_vector(8 downto 0);
      -- Read data output
      wb_fofb_processing_regs_ram_bank_9_data_o : out   std_logic_vector(31 downto 0);
      -- Read strobe input (active high)
      wb_fofb_processing_regs_ram_bank_9_rd_i : in    std_logic;
      -- Write data input
      wb_fofb_processing_regs_ram_bank_9_data_i : in    std_logic_vector(31 downto 0);
      -- Write strobe (active high)
      wb_fofb_processing_regs_ram_bank_9_wr_i : in    std_logic;
      -- Ports for RAM: FOFB PROCESSING RAM bank for register map
      wb_fofb_processing_regs_ram_bank_10_addr_i : in    std_logic_vector(8 downto 0);
      -- Read data output
      wb_fofb_processing_regs_ram_bank_10_data_o : out   std_logic_vector(31 downto 0);
      -- Read strobe input (active high)
      wb_fofb_processing_regs_ram_bank_10_rd_i : in    std_logic;
      -- Write data input
      wb_fofb_processing_regs_ram_bank_10_data_i : in    std_logic_vector(31 downto 0);
      -- Write strobe (active high)
      wb_fofb_processing_regs_ram_bank_10_wr_i : in    std_logic;
      -- Ports for RAM: FOFB PROCESSING RAM bank for register map
      wb_fofb_processing_regs_ram_bank_11_addr_i : in    std_logic_vector(8 downto 0);
      -- Read data output
      wb_fofb_processing_regs_ram_bank_11_data_o : out   std_logic_vector(31 downto 0);
      -- Read strobe input (active high)
      wb_fofb_processing_regs_ram_bank_11_rd_i : in    std_logic;
      -- Write data input
      wb_fofb_processing_regs_ram_bank_11_data_i : in    std_logic_vector(31 downto 0);
      -- Write strobe (active high)
      wb_fofb_processing_regs_ram_bank_11_wr_i : in    std_logic
    );
  end component wb_fofb_processing_regs;
end package dot_prod_pkg;
