package wb_fofb_processing_regs_consts_pkg is
  constant c_WB_FOFB_PROCESSING_REGS_SIZE : Natural := 53248;
  constant c_WB_FOFB_PROCESSING_REGS_FIXED_POINT_POS_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_FIXED_POINT_POS_SIZE : Natural := 64;
  constant c_WB_FOFB_PROCESSING_REGS_FIXED_POINT_POS_COEFF_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_FIXED_POINT_POS_COEFF_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_FIXED_POINT_POS_ACCS_GAINS_ADDR : Natural := 16#4#;
  constant c_WB_FOFB_PROCESSING_REGS_FIXED_POINT_POS_ACCS_GAINS_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_LOOP_INTLK_ADDR : Natural := 16#40#;
  constant c_WB_FOFB_PROCESSING_REGS_LOOP_INTLK_SIZE : Natural := 64;
  constant c_WB_FOFB_PROCESSING_REGS_LOOP_INTLK_CTL_ADDR : Natural := 16#40#;
  constant c_WB_FOFB_PROCESSING_REGS_LOOP_INTLK_CTL_STA_CLR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_LOOP_INTLK_CTL_SRC_EN_ORB_DISTORT_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_LOOP_INTLK_CTL_SRC_EN_PACKET_LOSS_OFFSET : Natural := 2;
  constant c_WB_FOFB_PROCESSING_REGS_LOOP_INTLK_STA_ADDR : Natural := 16#44#;
  constant c_WB_FOFB_PROCESSING_REGS_LOOP_INTLK_STA_ORB_DISTORT_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_LOOP_INTLK_STA_PACKET_LOSS_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_LOOP_INTLK_ORB_DISTORT_LIMIT_ADDR : Natural := 16#48#;
  constant c_WB_FOFB_PROCESSING_REGS_LOOP_INTLK_ORB_DISTORT_LIMIT_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_LOOP_INTLK_MIN_NUM_PKTS_ADDR : Natural := 16#4c#;
  constant c_WB_FOFB_PROCESSING_REGS_LOOP_INTLK_MIN_NUM_PKTS_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SP_DECIM_RATIO_MAX_ADDR : Natural := 16#80#;
  constant c_WB_FOFB_PROCESSING_REGS_SP_DECIM_RATIO_MAX_CTE_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_SPS_RAM_BANK_ADDR : Natural := 16#800#;
  constant c_WB_FOFB_PROCESSING_REGS_SPS_RAM_BANK_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_SPS_RAM_BANK_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_ADDR : Natural := 16#1000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_SIZE : Natural := 49152;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_ADDR : Natural := 16#1000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_SIZE : Natural := 4096;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_COEFF_RAM_BANK_ADDR : Natural := 16#1000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_COEFF_RAM_BANK_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_COEFF_RAM_BANK_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_ACC_ADDR : Natural := 16#1800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_ACC_SIZE : Natural := 32;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_ACC_CTL_ADDR : Natural := 16#1800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_ACC_CTL_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_ACC_CTL_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_ACC_GAIN_ADDR : Natural := 16#1804#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_ACC_GAIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_SP_LIMITS_ADDR : Natural := 16#1820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_SP_LIMITS_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_SP_LIMITS_MAX_ADDR : Natural := 16#1820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_SP_LIMITS_MAX_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_SP_LIMITS_MIN_ADDR : Natural := 16#1824#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_SP_LIMITS_MIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_SP_DECIM_ADDR : Natural := 16#1828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_SP_DECIM_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_SP_DECIM_DATA_ADDR : Natural := 16#1828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_SP_DECIM_DATA_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_SP_DECIM_RATIO_ADDR : Natural := 16#182c#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_0_SP_DECIM_RATIO_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_ADDR : Natural := 16#2000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_SIZE : Natural := 4096;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_COEFF_RAM_BANK_ADDR : Natural := 16#2000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_COEFF_RAM_BANK_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_COEFF_RAM_BANK_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_ACC_ADDR : Natural := 16#2800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_ACC_SIZE : Natural := 32;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_ACC_CTL_ADDR : Natural := 16#2800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_ACC_CTL_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_ACC_CTL_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_ACC_GAIN_ADDR : Natural := 16#2804#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_ACC_GAIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_SP_LIMITS_ADDR : Natural := 16#2820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_SP_LIMITS_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_SP_LIMITS_MAX_ADDR : Natural := 16#2820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_SP_LIMITS_MAX_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_SP_LIMITS_MIN_ADDR : Natural := 16#2824#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_SP_LIMITS_MIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_SP_DECIM_ADDR : Natural := 16#2828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_SP_DECIM_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_SP_DECIM_DATA_ADDR : Natural := 16#2828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_SP_DECIM_DATA_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_SP_DECIM_RATIO_ADDR : Natural := 16#282c#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_1_SP_DECIM_RATIO_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_ADDR : Natural := 16#3000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_SIZE : Natural := 4096;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_COEFF_RAM_BANK_ADDR : Natural := 16#3000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_COEFF_RAM_BANK_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_COEFF_RAM_BANK_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_ACC_ADDR : Natural := 16#3800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_ACC_SIZE : Natural := 32;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_ACC_CTL_ADDR : Natural := 16#3800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_ACC_CTL_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_ACC_CTL_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_ACC_GAIN_ADDR : Natural := 16#3804#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_ACC_GAIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_SP_LIMITS_ADDR : Natural := 16#3820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_SP_LIMITS_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_SP_LIMITS_MAX_ADDR : Natural := 16#3820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_SP_LIMITS_MAX_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_SP_LIMITS_MIN_ADDR : Natural := 16#3824#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_SP_LIMITS_MIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_SP_DECIM_ADDR : Natural := 16#3828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_SP_DECIM_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_SP_DECIM_DATA_ADDR : Natural := 16#3828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_SP_DECIM_DATA_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_SP_DECIM_RATIO_ADDR : Natural := 16#382c#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_2_SP_DECIM_RATIO_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_ADDR : Natural := 16#4000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_SIZE : Natural := 4096;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_COEFF_RAM_BANK_ADDR : Natural := 16#4000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_COEFF_RAM_BANK_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_COEFF_RAM_BANK_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_ACC_ADDR : Natural := 16#4800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_ACC_SIZE : Natural := 32;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_ACC_CTL_ADDR : Natural := 16#4800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_ACC_CTL_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_ACC_CTL_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_ACC_GAIN_ADDR : Natural := 16#4804#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_ACC_GAIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_SP_LIMITS_ADDR : Natural := 16#4820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_SP_LIMITS_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_SP_LIMITS_MAX_ADDR : Natural := 16#4820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_SP_LIMITS_MAX_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_SP_LIMITS_MIN_ADDR : Natural := 16#4824#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_SP_LIMITS_MIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_SP_DECIM_ADDR : Natural := 16#4828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_SP_DECIM_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_SP_DECIM_DATA_ADDR : Natural := 16#4828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_SP_DECIM_DATA_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_SP_DECIM_RATIO_ADDR : Natural := 16#482c#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_3_SP_DECIM_RATIO_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_ADDR : Natural := 16#5000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_SIZE : Natural := 4096;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_COEFF_RAM_BANK_ADDR : Natural := 16#5000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_COEFF_RAM_BANK_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_COEFF_RAM_BANK_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_ACC_ADDR : Natural := 16#5800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_ACC_SIZE : Natural := 32;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_ACC_CTL_ADDR : Natural := 16#5800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_ACC_CTL_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_ACC_CTL_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_ACC_GAIN_ADDR : Natural := 16#5804#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_ACC_GAIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_SP_LIMITS_ADDR : Natural := 16#5820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_SP_LIMITS_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_SP_LIMITS_MAX_ADDR : Natural := 16#5820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_SP_LIMITS_MAX_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_SP_LIMITS_MIN_ADDR : Natural := 16#5824#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_SP_LIMITS_MIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_SP_DECIM_ADDR : Natural := 16#5828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_SP_DECIM_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_SP_DECIM_DATA_ADDR : Natural := 16#5828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_SP_DECIM_DATA_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_SP_DECIM_RATIO_ADDR : Natural := 16#582c#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_4_SP_DECIM_RATIO_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_ADDR : Natural := 16#6000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_SIZE : Natural := 4096;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_COEFF_RAM_BANK_ADDR : Natural := 16#6000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_COEFF_RAM_BANK_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_COEFF_RAM_BANK_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_ACC_ADDR : Natural := 16#6800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_ACC_SIZE : Natural := 32;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_ACC_CTL_ADDR : Natural := 16#6800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_ACC_CTL_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_ACC_CTL_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_ACC_GAIN_ADDR : Natural := 16#6804#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_ACC_GAIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_SP_LIMITS_ADDR : Natural := 16#6820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_SP_LIMITS_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_SP_LIMITS_MAX_ADDR : Natural := 16#6820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_SP_LIMITS_MAX_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_SP_LIMITS_MIN_ADDR : Natural := 16#6824#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_SP_LIMITS_MIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_SP_DECIM_ADDR : Natural := 16#6828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_SP_DECIM_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_SP_DECIM_DATA_ADDR : Natural := 16#6828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_SP_DECIM_DATA_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_SP_DECIM_RATIO_ADDR : Natural := 16#682c#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_5_SP_DECIM_RATIO_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_ADDR : Natural := 16#7000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_SIZE : Natural := 4096;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_COEFF_RAM_BANK_ADDR : Natural := 16#7000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_COEFF_RAM_BANK_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_COEFF_RAM_BANK_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_ACC_ADDR : Natural := 16#7800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_ACC_SIZE : Natural := 32;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_ACC_CTL_ADDR : Natural := 16#7800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_ACC_CTL_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_ACC_CTL_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_ACC_GAIN_ADDR : Natural := 16#7804#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_ACC_GAIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_SP_LIMITS_ADDR : Natural := 16#7820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_SP_LIMITS_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_SP_LIMITS_MAX_ADDR : Natural := 16#7820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_SP_LIMITS_MAX_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_SP_LIMITS_MIN_ADDR : Natural := 16#7824#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_SP_LIMITS_MIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_SP_DECIM_ADDR : Natural := 16#7828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_SP_DECIM_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_SP_DECIM_DATA_ADDR : Natural := 16#7828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_SP_DECIM_DATA_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_SP_DECIM_RATIO_ADDR : Natural := 16#782c#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_6_SP_DECIM_RATIO_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_ADDR : Natural := 16#8000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_SIZE : Natural := 4096;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_COEFF_RAM_BANK_ADDR : Natural := 16#8000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_COEFF_RAM_BANK_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_COEFF_RAM_BANK_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_ACC_ADDR : Natural := 16#8800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_ACC_SIZE : Natural := 32;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_ACC_CTL_ADDR : Natural := 16#8800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_ACC_CTL_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_ACC_CTL_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_ACC_GAIN_ADDR : Natural := 16#8804#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_ACC_GAIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_SP_LIMITS_ADDR : Natural := 16#8820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_SP_LIMITS_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_SP_LIMITS_MAX_ADDR : Natural := 16#8820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_SP_LIMITS_MAX_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_SP_LIMITS_MIN_ADDR : Natural := 16#8824#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_SP_LIMITS_MIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_SP_DECIM_ADDR : Natural := 16#8828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_SP_DECIM_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_SP_DECIM_DATA_ADDR : Natural := 16#8828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_SP_DECIM_DATA_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_SP_DECIM_RATIO_ADDR : Natural := 16#882c#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_7_SP_DECIM_RATIO_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_ADDR : Natural := 16#9000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_SIZE : Natural := 4096;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_COEFF_RAM_BANK_ADDR : Natural := 16#9000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_COEFF_RAM_BANK_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_COEFF_RAM_BANK_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_ACC_ADDR : Natural := 16#9800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_ACC_SIZE : Natural := 32;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_ACC_CTL_ADDR : Natural := 16#9800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_ACC_CTL_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_ACC_CTL_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_ACC_GAIN_ADDR : Natural := 16#9804#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_ACC_GAIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_SP_LIMITS_ADDR : Natural := 16#9820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_SP_LIMITS_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_SP_LIMITS_MAX_ADDR : Natural := 16#9820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_SP_LIMITS_MAX_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_SP_LIMITS_MIN_ADDR : Natural := 16#9824#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_SP_LIMITS_MIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_SP_DECIM_ADDR : Natural := 16#9828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_SP_DECIM_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_SP_DECIM_DATA_ADDR : Natural := 16#9828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_SP_DECIM_DATA_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_SP_DECIM_RATIO_ADDR : Natural := 16#982c#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_8_SP_DECIM_RATIO_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_ADDR : Natural := 16#a000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_SIZE : Natural := 4096;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_COEFF_RAM_BANK_ADDR : Natural := 16#a000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_COEFF_RAM_BANK_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_COEFF_RAM_BANK_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_ACC_ADDR : Natural := 16#a800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_ACC_SIZE : Natural := 32;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_ACC_CTL_ADDR : Natural := 16#a800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_ACC_CTL_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_ACC_CTL_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_ACC_GAIN_ADDR : Natural := 16#a804#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_ACC_GAIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_SP_LIMITS_ADDR : Natural := 16#a820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_SP_LIMITS_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_SP_LIMITS_MAX_ADDR : Natural := 16#a820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_SP_LIMITS_MAX_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_SP_LIMITS_MIN_ADDR : Natural := 16#a824#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_SP_LIMITS_MIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_SP_DECIM_ADDR : Natural := 16#a828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_SP_DECIM_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_SP_DECIM_DATA_ADDR : Natural := 16#a828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_SP_DECIM_DATA_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_SP_DECIM_RATIO_ADDR : Natural := 16#a82c#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_9_SP_DECIM_RATIO_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_ADDR : Natural := 16#b000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_SIZE : Natural := 4096;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_COEFF_RAM_BANK_ADDR : Natural := 16#b000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_COEFF_RAM_BANK_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_COEFF_RAM_BANK_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_ACC_ADDR : Natural := 16#b800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_ACC_SIZE : Natural := 32;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_ACC_CTL_ADDR : Natural := 16#b800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_ACC_CTL_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_ACC_CTL_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_ACC_GAIN_ADDR : Natural := 16#b804#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_ACC_GAIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_SP_LIMITS_ADDR : Natural := 16#b820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_SP_LIMITS_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_SP_LIMITS_MAX_ADDR : Natural := 16#b820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_SP_LIMITS_MAX_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_SP_LIMITS_MIN_ADDR : Natural := 16#b824#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_SP_LIMITS_MIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_SP_DECIM_ADDR : Natural := 16#b828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_SP_DECIM_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_SP_DECIM_DATA_ADDR : Natural := 16#b828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_SP_DECIM_DATA_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_SP_DECIM_RATIO_ADDR : Natural := 16#b82c#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_10_SP_DECIM_RATIO_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_ADDR : Natural := 16#c000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_SIZE : Natural := 4096;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_COEFF_RAM_BANK_ADDR : Natural := 16#c000#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_COEFF_RAM_BANK_SIZE : Natural := 4;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_COEFF_RAM_BANK_DATA_ADDR : Natural := 16#0#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_ACC_ADDR : Natural := 16#c800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_ACC_SIZE : Natural := 32;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_ACC_CTL_ADDR : Natural := 16#c800#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_ACC_CTL_CLEAR_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_ACC_CTL_FREEZE_OFFSET : Natural := 1;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_ACC_GAIN_ADDR : Natural := 16#c804#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_ACC_GAIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_SP_LIMITS_ADDR : Natural := 16#c820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_SP_LIMITS_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_SP_LIMITS_MAX_ADDR : Natural := 16#c820#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_SP_LIMITS_MAX_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_SP_LIMITS_MIN_ADDR : Natural := 16#c824#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_SP_LIMITS_MIN_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_SP_DECIM_ADDR : Natural := 16#c828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_SP_DECIM_SIZE : Natural := 8;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_SP_DECIM_DATA_ADDR : Natural := 16#c828#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_SP_DECIM_DATA_VAL_OFFSET : Natural := 0;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_SP_DECIM_RATIO_ADDR : Natural := 16#c82c#;
  constant c_WB_FOFB_PROCESSING_REGS_CH_11_SP_DECIM_RATIO_VAL_OFFSET : Natural := 0;
end package wb_fofb_processing_regs_consts_pkg;
